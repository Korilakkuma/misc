module m_fpga();
endmodule
